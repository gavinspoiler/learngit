module github_test();
endmodule